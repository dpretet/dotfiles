`timescale 1 ns / 1 ps
`default_nettype none

module ModuleName

    #(
    parameter NAME = 0
    )(
    input         aclk,
    input         aresetn,
    input         wen,
    input  [15:0] wdata,
    output logic  wout
    );


endmodule

`resetall
