`timescale 1 ns / 1 ps
`default_nettype none

module ModuleName

    #(
    parameter NAME = 0
    )(
    input  wire aclk,
    input  wire arstn,
    output wire out
    );

endmodule

`resetall
